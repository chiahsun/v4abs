module top(clk);

initial begin
    a.sub.b.in1 = 1'b1;
end

endmodule
