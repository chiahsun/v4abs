module A(reset);

parameter A = 10;
endmodule
