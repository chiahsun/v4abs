always @ (*) begin
    next_state = state;
    next_reg_i = reg_i;
end
