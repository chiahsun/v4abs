`timescale 10ns/1ns

`include "./sram_1024x8_t13.v"

module sram_ctrl(clk, reset, sram_in_ctrl, sram_in, sram_out);

input        clk;
input        reset;
input  [1:0] sram_in_ctrl;
input  [7:0] sram_in;
output [7:0] sram_out;



reg   [9:0] sram_write_addr;
wire   [9:0] sram_read_addr;
wire  [9:0] sram_addr;
wire  [7:0] tmp;

reg sram_en, sram_w_r;
reg [7:0] internal_counter;

reg    [7:0] sram_data_in;
reg    [7:0] sram_data_out;
reg sram_CEB;
always @ (posedge clk) begin
    sram_data_in  <= (reset) ? 0 : sram_in;
    sram_data_out <= (reset) ? 0 : tmp;
    sram_en       <= (reset) ? 0 : sram_in_ctrl[1];
    sram_w_r      <= (reset) ? 0 : sram_in_ctrl[0];
end

assign sram_addr = (sram_w_r) ? sram_write_addr : sram_read_addr;
assign sram_read_addr = sram_write_addr -128 + internal_counter;
reg [7:0] cnt;
wire [7:0] dbg_cnt;
assign dbg_cnt = cnt;
always @ (posedge clk) begin
    if(!sram_en) cnt <= 0;
    else cnt <= (cnt == 8'h82) ? 0 : cnt+1'b1;
end
always @ (posedge clk) begin
    if(!sram_en) internal_counter <= 0;
    else
         if(!sram_w_r) 
            internal_counter <= (cnt == 8'h82) 
                             ? 0
                             : internal_counter + 1'b1;
end
always @ (posedge clk) begin
    if(reset) begin
        sram_CEB <= 1'b1;
        sram_write_addr <= 0;
    end
    else begin 
        sram_CEB <= 1'b0;
        if(sram_en && sram_w_r) 
            sram_write_addr <= sram_write_addr + 1'b1 ;
    end
end


sram_1024x8_t13 my_ram(.A(sram_addr),
                   .D(sram_data_in),
                   .CLK(~clk),
                   .CEN(sram_CEB),
                   .WEN(~sram_w_r),
                   .Q(tmp) );
assign sram_out = tmp;

endmodule
module comparator(d1_in, d2_in, d1_out, d2_out);
    input  [7:0] d1_in, d2_in;
    output [7:0] d1_out, d2_out;
    assign {d2_out,d1_out} = (d1_in > d2_in) ? {d1_in,d2_in} : {d2_in,d1_in};
endmodule


module bsort(data_in, data_out);


input   [511:0] data_in;
output  [511:0] data_out;

wire[7:0] a10v1, a10v10, a10v11, a10v12, a10v13, a10v14, a10v15, a10v16, a10v17, a10v18,     
a10v19, a10v2, a10v20, a10v21, a10v22, a10v23, a10v24, a10v25, a10v26, a10v27,     
a10v28, a10v29, a10v3, a10v30, a10v31, a10v32, a10v33, a10v34, a10v35, a10v36,     
a10v37, a10v38, a10v39, a10v4, a10v40, a10v41, a10v42, a10v43, a10v44, a10v45,     
a10v46, a10v47, a10v48, a10v49, a10v5, a10v50, a10v51, a10v52, a10v53, a10v54,     
a10v55, a10v56, a10v57, a10v58, a10v59, a10v6, a10v60, a10v61, a10v62, a10v7,     
a10v8, a10v9, a11v1, a11v10, a11v11, a11v12, a11v13, a11v14, a11v15, a11v16,     
a11v17, a11v18, a11v19, a11v2, a11v20, a11v21, a11v22, a11v23, a11v24, a11v25,     
a11v26, a11v27, a11v28, a11v29, a11v3, a11v30, a11v31, a11v32, a11v33, a11v34,     
a11v35, a11v36, a11v37, a11v38, a11v39, a11v4, a11v40, a11v41, a11v42, a11v43,     
a11v44, a11v45, a11v46, a11v47, a11v48, a11v49, a11v5, a11v50, a11v51, a11v52,     
a11v53, a11v54, a11v55, a11v56, a11v57, a11v58, a11v59, a11v6, a11v60, a11v61,     
a11v62, a11v7, a11v8, a11v9, a12v1, a12v10, a12v11, a12v12, a12v13, a12v14,     
a12v15, a12v16, a12v17, a12v18, a12v19, a12v2, a12v20, a12v21, a12v22, a12v23,     
a12v24, a12v25, a12v26, a12v27, a12v28, a12v29, a12v3, a12v30, a12v31, a12v32,     
a12v33, a12v34, a12v35, a12v36, a12v37, a12v38, a12v39, a12v4, a12v40, a12v41,     
a12v42, a12v43, a12v44, a12v45, a12v46, a12v47, a12v48, a12v49, a12v5, a12v50,     
a12v51, a12v52, a12v53, a12v54, a12v55, a12v56, a12v57, a12v58, a12v59, a12v6,     
a12v60, a12v61, a12v62, a12v7, a12v8, a12v9, a13v10, a13v11, a13v12, a13v13,     
a13v14, a13v15, a13v16, a13v17, a13v18, a13v19, a13v2, a13v20, a13v21, a13v22,     
a13v23, a13v24, a13v25, a13v26, a13v27, a13v28, a13v29, a13v3, a13v30, a13v33,     
a13v34, a13v35, a13v36, a13v37, a13v38, a13v39, a13v4, a13v40, a13v41, a13v42,     
a13v43, a13v44, a13v45, a13v46, a13v47, a13v48, a13v49, a13v5, a13v50, a13v51,     
a13v52, a13v53, a13v54, a13v55, a13v56, a13v57, a13v58, a13v59, a13v6, a13v60,     
a13v61, a13v7, a13v8, a13v9, a14v10, a14v11, a14v12, a14v13, a14v14, a14v15,     
a14v16, a14v17, a14v18, a14v19, a14v2, a14v20, a14v21, a14v22, a14v23, a14v24,     
a14v25, a14v26, a14v27, a14v28, a14v29, a14v3, a14v30, a14v33, a14v34, a14v35,     
a14v36, a14v37, a14v38, a14v39, a14v4, a14v40, a14v41, a14v42, a14v43, a14v44,     
a14v45, a14v46, a14v47, a14v48, a14v49, a14v5, a14v50, a14v51, a14v52, a14v53,     
a14v54, a14v55, a14v56, a14v57, a14v58, a14v59, a14v6, a14v60, a14v61, a14v7,     
a14v8, a14v9, a15v10, a15v11, a15v12, a15v13, a15v14, a15v15, a15v16, a15v17,     
a15v18, a15v19, a15v2, a15v20, a15v21, a15v22, a15v23, a15v24, a15v25, a15v26,     
a15v27, a15v28, a15v29, a15v3, a15v30, a15v33, a15v34, a15v35, a15v36, a15v37,     
a15v38, a15v39, a15v4, a15v40, a15v41, a15v42, a15v43, a15v44, a15v45, a15v46,     
a15v47, a15v48, a15v49, a15v5, a15v50, a15v51, a15v52, a15v53, a15v54, a15v55,     
a15v56, a15v57, a15v58, a15v59, a15v6, a15v60, a15v61, a15v7, a15v8, a15v9,     
a16v10, a16v11, a16v12, a16v13, a16v14, a16v16, a16v17, a16v18, a16v19, a16v2,     
a16v20, a16v21, a16v22, a16v23, a16v24, a16v25, a16v26, a16v27, a16v28, a16v29,     
a16v30, a16v33, a16v34, a16v35, a16v36, a16v37, a16v38, a16v39, a16v4, a16v40,     
a16v41, a16v42, a16v43, a16v44, a16v45, a16v46, a16v47, a16v49, a16v5, a16v50,     
a16v51, a16v52, a16v53, a16v54, a16v55, a16v56, a16v57, a16v58, a16v59, a16v6,     
a16v61, a16v7, a16v8, a16v9, a17v10, a17v11, a17v12, a17v13, a17v14, a17v17,     
a17v18, a17v19, a17v20, a17v21, a17v22, a17v23, a17v24, a17v25, a17v26, a17v27,     
a17v28, a17v29, a17v34, a17v35, a17v36, a17v37, a17v38, a17v39, a17v4, a17v40,     
a17v41, a17v42, a17v43, a17v44, a17v45, a17v46, a17v49, a17v5, a17v50, a17v51,     
a17v52, a17v53, a17v54, a17v55, a17v57, a17v58, a17v59, a17v6, a17v8, a17v9,     
a18v10, a18v11, a18v12, a18v13, a18v14, a18v17, a18v18, a18v19, a18v20, a18v21,     
a18v22, a18v23, a18v24, a18v25, a18v26, a18v27, a18v28, a18v29, a18v34, a18v35,     
a18v36, a18v37, a18v38, a18v39, a18v4, a18v40, a18v41, a18v42, a18v43, a18v44,     
a18v45, a18v46, a18v49, a18v5, a18v50, a18v51, a18v52, a18v53, a18v54, a18v55,     
a18v57, a18v58, a18v59, a18v6, a18v8, a18v9, a19v10, a19v11, a19v12, a19v13,     
a19v17, a19v18, a19v19, a19v20, a19v21, a19v22, a19v23, a19v25, a19v26, a19v27,     
a19v29, a19v34, a19v36, a19v37, a19v38, a19v40, a19v41, a19v42, a19v43, a19v44,     
a19v45, a19v46, a19v5, a19v50, a19v51, a19v52, a19v53, a19v54, a19v58, a19v9,     
a1v0, a1v1, a1v10, a1v11, a1v12, a1v13, a1v14, a1v15, a1v16, a1v17,     
a1v18, a1v19, a1v2, a1v20, a1v21, a1v22, a1v23, a1v24, a1v25, a1v26,     
a1v27, a1v28, a1v29, a1v3, a1v30, a1v31, a1v32, a1v33, a1v34, a1v35,     
a1v36, a1v37, a1v38, a1v39, a1v4, a1v40, a1v41, a1v42, a1v43, a1v44,     
a1v45, a1v46, a1v47, a1v48, a1v49, a1v5, a1v50, a1v51, a1v52, a1v53,     
a1v54, a1v55, a1v56, a1v57, a1v58, a1v59, a1v6, a1v60, a1v61, a1v62,     
a1v63, a1v7, a1v8, a1v9, a20v10, a20v11, a20v13, a20v18, a20v19, a20v20,     
a20v21, a20v22, a20v25, a20v26, a20v27, a20v36, a20v37, a20v38, a20v41, a20v42,     
a20v43, a20v44, a20v45, a20v50, a20v52, a20v53, a20v54, a20v9, a21v10, a21v18,     
a21v20, a21v21, a21v22, a21v26, a21v37, a21v41, a21v42, a21v43, a21v45, a21v53,     
a22v21, a22v42, a2v0, a2v1, a2v10, a2v11, a2v12, a2v13, a2v14, a2v15,     
a2v16, a2v17, a2v18, a2v19, a2v2, a2v20, a2v21, a2v22, a2v23, a2v24,     
a2v25, a2v26, a2v27, a2v28, a2v29, a2v3, a2v30, a2v31, a2v32, a2v33,     
a2v34, a2v35, a2v36, a2v37, a2v38, a2v39, a2v4, a2v40, a2v41, a2v42,     
a2v43, a2v44, a2v45, a2v46, a2v47, a2v48, a2v49, a2v5, a2v50, a2v51,     
a2v52, a2v53, a2v54, a2v55, a2v56, a2v57, a2v58, a2v59, a2v6, a2v60,     
a2v61, a2v62, a2v63, a2v7, a2v8, a2v9, a3v0, a3v1, a3v10, a3v11,     
a3v12, a3v13, a3v14, a3v15, a3v16, a3v17, a3v18, a3v19, a3v2, a3v20,     
a3v21, a3v22, a3v23, a3v24, a3v25, a3v26, a3v27, a3v28, a3v29, a3v3,     
a3v30, a3v31, a3v32, a3v33, a3v34, a3v35, a3v36, a3v37, a3v38, a3v39,     
a3v4, a3v40, a3v41, a3v42, a3v43, a3v44, a3v45, a3v46, a3v47, a3v48,     
a3v49, a3v5, a3v50, a3v51, a3v52, a3v53, a3v54, a3v55, a3v56, a3v57,     
a3v58, a3v59, a3v6, a3v60, a3v61, a3v62, a3v63, a3v7, a3v8, a3v9,     
a4v0, a4v1, a4v10, a4v11, a4v12, a4v13, a4v14, a4v15, a4v16, a4v17,     
a4v18, a4v19, a4v2, a4v20, a4v21, a4v22, a4v23, a4v24, a4v25, a4v26,     
a4v27, a4v28, a4v29, a4v3, a4v30, a4v31, a4v32, a4v33, a4v34, a4v35,     
a4v36, a4v37, a4v38, a4v39, a4v4, a4v40, a4v41, a4v42, a4v43, a4v44,     
a4v45, a4v46, a4v47, a4v48, a4v49, a4v5, a4v50, a4v51, a4v52, a4v53,     
a4v54, a4v55, a4v56, a4v57, a4v58, a4v59, a4v6, a4v60, a4v61, a4v62,     
a4v63, a4v7, a4v8, a4v9, a5v0, a5v1, a5v10, a5v11, a5v12, a5v13,     
a5v14, a5v15, a5v16, a5v17, a5v18, a5v19, a5v2, a5v20, a5v21, a5v22,     
a5v23, a5v24, a5v25, a5v26, a5v27, a5v28, a5v29, a5v3, a5v30, a5v31,     
a5v32, a5v33, a5v34, a5v35, a5v36, a5v37, a5v38, a5v39, a5v4, a5v40,     
a5v41, a5v42, a5v43, a5v44, a5v45, a5v46, a5v47, a5v48, a5v49, a5v5,     
a5v50, a5v51, a5v52, a5v53, a5v54, a5v55, a5v56, a5v57, a5v58, a5v59,     
a5v6, a5v60, a5v61, a5v62, a5v63, a5v7, a5v8, a5v9, a6v0, a6v1,     
a6v10, a6v11, a6v12, a6v13, a6v14, a6v15, a6v16, a6v17, a6v18, a6v19,     
a6v2, a6v20, a6v21, a6v22, a6v23, a6v24, a6v25, a6v26, a6v27, a6v28,     
a6v29, a6v3, a6v30, a6v31, a6v32, a6v33, a6v34, a6v35, a6v36, a6v37,     
a6v38, a6v39, a6v4, a6v40, a6v41, a6v42, a6v43, a6v44, a6v45, a6v46,     
a6v47, a6v48, a6v49, a6v5, a6v50, a6v51, a6v52, a6v53, a6v54, a6v55,     
a6v56, a6v57, a6v58, a6v59, a6v6, a6v60, a6v61, a6v62, a6v63, a6v7,     
a6v8, a6v9, a7v0, a7v1, a7v10, a7v11, a7v12, a7v13, a7v14, a7v15,     
a7v16, a7v17, a7v18, a7v19, a7v2, a7v20, a7v21, a7v22, a7v23, a7v24,     
a7v25, a7v26, a7v27, a7v28, a7v29, a7v3, a7v30, a7v31, a7v32, a7v33,     
a7v34, a7v35, a7v36, a7v37, a7v38, a7v39, a7v4, a7v40, a7v41, a7v42,     
a7v43, a7v44, a7v45, a7v46, a7v47, a7v48, a7v49, a7v5, a7v50, a7v51,     
a7v52, a7v53, a7v54, a7v55, a7v56, a7v57, a7v58, a7v59, a7v6, a7v60,     
a7v61, a7v62, a7v63, a7v7, a7v8, a7v9, a8v1, a8v10, a8v11, a8v12,     
a8v13, a8v14, a8v15, a8v16, a8v17, a8v18, a8v19, a8v2, a8v20, a8v21,     
a8v22, a8v23, a8v24, a8v25, a8v26, a8v27, a8v28, a8v29, a8v3, a8v30,     
a8v31, a8v32, a8v33, a8v34, a8v35, a8v36, a8v37, a8v38, a8v39, a8v4,     
a8v40, a8v41, a8v42, a8v43, a8v44, a8v45, a8v46, a8v47, a8v48, a8v49,     
a8v5, a8v50, a8v51, a8v52, a8v53, a8v54, a8v55, a8v56, a8v57, a8v58,     
a8v59, a8v6, a8v60, a8v61, a8v62, a8v7, a8v8, a8v9, a9v1, a9v10,     
a9v11, a9v12, a9v13, a9v14, a9v15, a9v16, a9v17, a9v18, a9v19, a9v2,     
a9v20, a9v21, a9v22, a9v23, a9v24, a9v25, a9v26, a9v27, a9v28, a9v29,     
a9v3, a9v30, a9v31, a9v32, a9v33, a9v34, a9v35, a9v36, a9v37, a9v38,     
a9v39, a9v4, a9v40, a9v41, a9v42, a9v43, a9v44, a9v45, a9v46, a9v47,     
a9v48, a9v49, a9v5, a9v50, a9v51, a9v52, a9v53, a9v54, a9v55, a9v56,     
a9v57, a9v58, a9v59, a9v6, a9v60, a9v61, a9v62, a9v7, a9v8, a9v9    
;


assign a1v0 = data_in[7:0];
assign a1v1 = data_in[15:8];
assign a1v2 = data_in[23:16];
assign a1v3 = data_in[31:24];
assign a1v4 = data_in[39:32];
assign a1v5 = data_in[47:40];
assign a1v6 = data_in[55:48];
assign a1v7 = data_in[63:56];
assign a1v8 = data_in[71:64];
assign a1v9 = data_in[79:72];
assign a1v10 = data_in[87:80];
assign a1v11 = data_in[95:88];
assign a1v12 = data_in[103:96];
assign a1v13 = data_in[111:104];
assign a1v14 = data_in[119:112];
assign a1v15 = data_in[127:120];
assign a1v16 = data_in[135:128];
assign a1v17 = data_in[143:136];
assign a1v18 = data_in[151:144];
assign a1v19 = data_in[159:152];
assign a1v20 = data_in[167:160];
assign a1v21 = data_in[175:168];
assign a1v22 = data_in[183:176];
assign a1v23 = data_in[191:184];
assign a1v24 = data_in[199:192];
assign a1v25 = data_in[207:200];
assign a1v26 = data_in[215:208];
assign a1v27 = data_in[223:216];
assign a1v28 = data_in[231:224];
assign a1v29 = data_in[239:232];
assign a1v30 = data_in[247:240];
assign a1v31 = data_in[255:248];
assign a1v32 = data_in[263:256];
assign a1v33 = data_in[271:264];
assign a1v34 = data_in[279:272];
assign a1v35 = data_in[287:280];
assign a1v36 = data_in[295:288];
assign a1v37 = data_in[303:296];
assign a1v38 = data_in[311:304];
assign a1v39 = data_in[319:312];
assign a1v40 = data_in[327:320];
assign a1v41 = data_in[335:328];
assign a1v42 = data_in[343:336];
assign a1v43 = data_in[351:344];
assign a1v44 = data_in[359:352];
assign a1v45 = data_in[367:360];
assign a1v46 = data_in[375:368];
assign a1v47 = data_in[383:376];
assign a1v48 = data_in[391:384];
assign a1v49 = data_in[399:392];
assign a1v50 = data_in[407:400];
assign a1v51 = data_in[415:408];
assign a1v52 = data_in[423:416];
assign a1v53 = data_in[431:424];
assign a1v54 = data_in[439:432];
assign a1v55 = data_in[447:440];
assign a1v56 = data_in[455:448];
assign a1v57 = data_in[463:456];
assign a1v58 = data_in[471:464];
assign a1v59 = data_in[479:472];
assign a1v60 = data_in[487:480];
assign a1v61 = data_in[495:488];
assign a1v62 = data_in[503:496];
assign a1v63 = data_in[511:504];

assign data_out[7:0] = a7v0;
assign data_out[15:8] = a12v1;
assign data_out[23:16] = a16v2;
assign data_out[31:24] = a15v3;
assign data_out[39:32] = a18v4;
assign data_out[47:40] = a19v5;
assign data_out[55:48] = a18v6;
assign data_out[63:56] = a16v7;
assign data_out[71:64] = a18v8;
assign data_out[79:72] = a20v9;
assign data_out[87:80] = a21v10;
assign data_out[95:88] = a20v11;
assign data_out[103:96] = a19v12;
assign data_out[111:104] = a20v13;
assign data_out[119:112] = a18v14;
assign data_out[127:120] = a15v15;
assign data_out[135:128] = a16v16;
assign data_out[143:136] = a19v17;
assign data_out[151:144] = a21v18;
assign data_out[159:152] = a20v19;
assign data_out[167:160] = a21v20;
assign data_out[175:168] = a22v21;
assign data_out[183:176] = a21v22;
assign data_out[191:184] = a19v23;
assign data_out[199:192] = a18v24;
assign data_out[207:200] = a20v25;
assign data_out[215:208] = a21v26;
assign data_out[223:216] = a20v27;
assign data_out[231:224] = a18v28;
assign data_out[239:232] = a19v29;
assign data_out[247:240] = a16v30;
assign data_out[255:248] = a12v31;
assign data_out[263:256] = a12v32;
assign data_out[271:264] = a16v33;
assign data_out[279:272] = a19v34;
assign data_out[287:280] = a18v35;
assign data_out[295:288] = a20v36;
assign data_out[303:296] = a21v37;
assign data_out[311:304] = a20v38;
assign data_out[319:312] = a18v39;
assign data_out[327:320] = a19v40;
assign data_out[335:328] = a21v41;
assign data_out[343:336] = a22v42;
assign data_out[351:344] = a21v43;
assign data_out[359:352] = a20v44;
assign data_out[367:360] = a21v45;
assign data_out[375:368] = a19v46;
assign data_out[383:376] = a16v47;
assign data_out[391:384] = a15v48;
assign data_out[399:392] = a18v49;
assign data_out[407:400] = a20v50;
assign data_out[415:408] = a19v51;
assign data_out[423:416] = a20v52;
assign data_out[431:424] = a21v53;
assign data_out[439:432] = a20v54;
assign data_out[447:440] = a18v55;
assign data_out[455:448] = a16v56;
assign data_out[463:456] = a18v57;
assign data_out[471:464] = a19v58;
assign data_out[479:472] = a18v59;
assign data_out[487:480] = a15v60;
assign data_out[495:488] = a16v61;
assign data_out[503:496] = a12v62;
assign data_out[511:504] = a7v63;


comparator c0 (a1v0, a1v1, a2v0, a2v1);
comparator c1 (a1v2, a1v3, a2v2, a2v3);
comparator c2 (a2v0, a2v2, a3v0, a3v2);
comparator c3 (a2v1, a2v3, a3v1, a3v3);
comparator c4 (a3v1, a3v2, a4v1, a4v2);
comparator c5 (a1v4, a1v5, a2v4, a2v5);
comparator c6 (a1v6, a1v7, a2v6, a2v7);
comparator c7 (a2v4, a2v6, a3v4, a3v6);
comparator c8 (a2v5, a2v7, a3v5, a3v7);
comparator c9 (a3v5, a3v6, a4v5, a4v6);
comparator c10 (a3v0, a3v4, a4v0, a4v4);
comparator c11 (a4v2, a4v6, a5v2, a5v6);
comparator c12 (a5v2, a4v4, a6v2, a5v4);
comparator c13 (a4v1, a4v5, a5v1, a5v5);
comparator c14 (a3v3, a3v7, a4v3, a4v7);
comparator c15 (a4v3, a5v5, a5v3, a6v5);
comparator c16 (a5v1, a6v2, a6v1, a7v2);
comparator c17 (a5v3, a5v4, a6v3, a6v4);
comparator c18 (a6v5, a5v6, a7v5, a6v6);
comparator c19 (a1v8, a1v9, a2v8, a2v9);
comparator c20 (a1v10, a1v11, a2v10, a2v11);
comparator c21 (a2v8, a2v10, a3v8, a3v10);
comparator c22 (a2v9, a2v11, a3v9, a3v11);
comparator c23 (a3v9, a3v10, a4v9, a4v10);
comparator c24 (a1v12, a1v13, a2v12, a2v13);
comparator c25 (a1v14, a1v15, a2v14, a2v15);
comparator c26 (a2v12, a2v14, a3v12, a3v14);
comparator c27 (a2v13, a2v15, a3v13, a3v15);
comparator c28 (a3v13, a3v14, a4v13, a4v14);
comparator c29 (a3v8, a3v12, a4v8, a4v12);
comparator c30 (a4v10, a4v14, a5v10, a5v14);
comparator c31 (a5v10, a4v12, a6v10, a5v12);
comparator c32 (a4v9, a4v13, a5v9, a5v13);
comparator c33 (a3v11, a3v15, a4v11, a4v15);
comparator c34 (a4v11, a5v13, a5v11, a6v13);
comparator c35 (a5v9, a6v10, a6v9, a7v10);
comparator c36 (a5v11, a5v12, a6v11, a6v12);
comparator c37 (a6v13, a5v14, a7v13, a6v14);
comparator c38 (a4v0, a4v8, a5v0, a5v8);
comparator c39 (a6v4, a6v12, a7v4, a7v12);
comparator c40 (a7v4, a5v8, a8v4, a6v8);
comparator c41 (a7v2, a7v10, a8v2, a8v10);
comparator c42 (a6v6, a6v14, a7v6, a7v14);
comparator c43 (a7v6, a8v10, a8v6, a9v10);
comparator c44 (a8v2, a8v4, a9v2, a9v4);
comparator c45 (a8v6, a6v8, a9v6, a7v8);
comparator c46 (a9v10, a7v12, a10v10, a8v12);
comparator c47 (a6v1, a6v9, a7v1, a7v9);
comparator c48 (a7v5, a7v13, a8v5, a8v13);
comparator c49 (a8v5, a7v9, a9v5, a8v9);
comparator c50 (a6v3, a6v11, a7v3, a7v11);
comparator c51 (a4v7, a4v15, a5v7, a5v15);
comparator c52 (a5v7, a7v11, a6v7, a8v11);
comparator c53 (a7v3, a9v5, a8v3, a10v5);
comparator c54 (a6v7, a8v9, a7v7, a9v9);
comparator c55 (a8v11, a8v13, a9v11, a9v13);
comparator c56 (a7v1, a9v2, a8v1, a10v2);
comparator c57 (a8v3, a9v4, a9v3, a10v4);
comparator c58 (a10v5, a9v6, a11v5, a10v6);
comparator c59 (a7v7, a7v8, a8v7, a8v8);
comparator c60 (a9v9, a10v10, a10v9, a11v10);
comparator c61 (a9v11, a8v12, a10v11, a9v12);
comparator c62 (a9v13, a7v14, a10v13, a8v14);
comparator c63 (a1v16, a1v17, a2v16, a2v17);
comparator c64 (a1v18, a1v19, a2v18, a2v19);
comparator c65 (a2v16, a2v18, a3v16, a3v18);
comparator c66 (a2v17, a2v19, a3v17, a3v19);
comparator c67 (a3v17, a3v18, a4v17, a4v18);
comparator c68 (a1v20, a1v21, a2v20, a2v21);
comparator c69 (a1v22, a1v23, a2v22, a2v23);
comparator c70 (a2v20, a2v22, a3v20, a3v22);
comparator c71 (a2v21, a2v23, a3v21, a3v23);
comparator c72 (a3v21, a3v22, a4v21, a4v22);
comparator c73 (a3v16, a3v20, a4v16, a4v20);
comparator c74 (a4v18, a4v22, a5v18, a5v22);
comparator c75 (a5v18, a4v20, a6v18, a5v20);
comparator c76 (a4v17, a4v21, a5v17, a5v21);
comparator c77 (a3v19, a3v23, a4v19, a4v23);
comparator c78 (a4v19, a5v21, a5v19, a6v21);
comparator c79 (a5v17, a6v18, a6v17, a7v18);
comparator c80 (a5v19, a5v20, a6v19, a6v20);
comparator c81 (a6v21, a5v22, a7v21, a6v22);
comparator c82 (a1v24, a1v25, a2v24, a2v25);
comparator c83 (a1v26, a1v27, a2v26, a2v27);
comparator c84 (a2v24, a2v26, a3v24, a3v26);
comparator c85 (a2v25, a2v27, a3v25, a3v27);
comparator c86 (a3v25, a3v26, a4v25, a4v26);
comparator c87 (a1v28, a1v29, a2v28, a2v29);
comparator c88 (a1v30, a1v31, a2v30, a2v31);
comparator c89 (a2v28, a2v30, a3v28, a3v30);
comparator c90 (a2v29, a2v31, a3v29, a3v31);
comparator c91 (a3v29, a3v30, a4v29, a4v30);
comparator c92 (a3v24, a3v28, a4v24, a4v28);
comparator c93 (a4v26, a4v30, a5v26, a5v30);
comparator c94 (a5v26, a4v28, a6v26, a5v28);
comparator c95 (a4v25, a4v29, a5v25, a5v29);
comparator c96 (a3v27, a3v31, a4v27, a4v31);
comparator c97 (a4v27, a5v29, a5v27, a6v29);
comparator c98 (a5v25, a6v26, a6v25, a7v26);
comparator c99 (a5v27, a5v28, a6v27, a6v28);
comparator c100 (a6v29, a5v30, a7v29, a6v30);
comparator c101 (a4v16, a4v24, a5v16, a5v24);
comparator c102 (a6v20, a6v28, a7v20, a7v28);
comparator c103 (a7v20, a5v24, a8v20, a6v24);
comparator c104 (a7v18, a7v26, a8v18, a8v26);
comparator c105 (a6v22, a6v30, a7v22, a7v30);
comparator c106 (a7v22, a8v26, a8v22, a9v26);
comparator c107 (a8v18, a8v20, a9v18, a9v20);
comparator c108 (a8v22, a6v24, a9v22, a7v24);
comparator c109 (a9v26, a7v28, a10v26, a8v28);
comparator c110 (a6v17, a6v25, a7v17, a7v25);
comparator c111 (a7v21, a7v29, a8v21, a8v29);
comparator c112 (a8v21, a7v25, a9v21, a8v25);
comparator c113 (a6v19, a6v27, a7v19, a7v27);
comparator c114 (a4v23, a4v31, a5v23, a5v31);
comparator c115 (a5v23, a7v27, a6v23, a8v27);
comparator c116 (a7v19, a9v21, a8v19, a10v21);
comparator c117 (a6v23, a8v25, a7v23, a9v25);
comparator c118 (a8v27, a8v29, a9v27, a9v29);
comparator c119 (a7v17, a9v18, a8v17, a10v18);
comparator c120 (a8v19, a9v20, a9v19, a10v20);
comparator c121 (a10v21, a9v22, a11v21, a10v22);
comparator c122 (a7v23, a7v24, a8v23, a8v24);
comparator c123 (a9v25, a10v26, a10v25, a11v26);
comparator c124 (a9v27, a8v28, a10v27, a9v28);
comparator c125 (a9v29, a7v30, a10v29, a8v30);
comparator c126 (a5v0, a5v16, a6v0, a6v16);
comparator c127 (a8v8, a8v24, a9v8, a9v24);
comparator c128 (a9v8, a6v16, a10v8, a7v16);
comparator c129 (a10v4, a10v20, a11v4, a11v20);
comparator c130 (a9v12, a9v28, a10v12, a10v28);
comparator c131 (a10v12, a11v20, a11v12, a12v20);
comparator c132 (a11v4, a10v8, a12v4, a11v8);
comparator c133 (a11v12, a7v16, a12v12, a8v16);
comparator c134 (a12v20, a9v24, a13v20, a10v24);
comparator c135 (a10v2, a10v18, a11v2, a11v18);
comparator c136 (a11v10, a11v26, a12v10, a12v26);
comparator c137 (a12v10, a11v18, a13v10, a12v18);
comparator c138 (a10v6, a10v22, a11v6, a11v22);
comparator c139 (a8v14, a8v30, a9v14, a9v30);
comparator c140 (a9v14, a11v22, a10v14, a12v22);
comparator c141 (a11v6, a13v10, a12v6, a14v10);
comparator c142 (a10v14, a12v18, a11v14, a13v18);
comparator c143 (a12v22, a12v26, a13v22, a13v26);
comparator c144 (a11v2, a12v4, a12v2, a13v4);
comparator c145 (a12v6, a11v8, a13v6, a12v8);
comparator c146 (a14v10, a12v12, a15v10, a13v12);
comparator c147 (a11v14, a8v16, a12v14, a9v16);
comparator c148 (a13v18, a13v20, a14v18, a14v20);
comparator c149 (a13v22, a10v24, a14v22, a11v24);
comparator c150 (a13v26, a10v28, a14v26, a11v28);
comparator c151 (a8v1, a8v17, a9v1, a9v17);
comparator c152 (a10v9, a10v25, a11v9, a11v25);
comparator c153 (a11v9, a9v17, a12v9, a10v17);
comparator c154 (a11v5, a11v21, a12v5, a12v21);
comparator c155 (a10v13, a10v29, a11v13, a11v29);
comparator c156 (a11v13, a12v21, a12v13, a13v21);
comparator c157 (a12v5, a12v9, a13v5, a13v9);
comparator c158 (a12v13, a10v17, a13v13, a11v17);
comparator c159 (a13v21, a11v25, a14v21, a12v25);
comparator c160 (a9v3, a9v19, a10v3, a10v19);
comparator c161 (a10v11, a10v27, a11v11, a11v27);
comparator c162 (a11v11, a10v19, a12v11, a11v19);
comparator c163 (a8v7, a8v23, a9v7, a9v23);
comparator c164 (a5v15, a5v31, a6v15, a6v31);
comparator c165 (a6v15, a9v23, a7v15, a10v23);
comparator c166 (a9v7, a12v11, a10v7, a13v11);
comparator c167 (a7v15, a11v19, a8v15, a12v19);
comparator c168 (a10v23, a11v27, a11v23, a12v27);
comparator c169 (a10v3, a13v5, a11v3, a14v5);
comparator c170 (a10v7, a13v9, a11v7, a14v9);
comparator c171 (a13v11, a13v13, a14v11, a14v13);
comparator c172 (a8v15, a11v17, a9v15, a12v17);
comparator c173 (a12v19, a14v21, a13v19, a15v21);
comparator c174 (a11v23, a12v25, a12v23, a13v25);
comparator c175 (a12v27, a11v29, a13v27, a12v29);
comparator c176 (a9v1, a12v2, a10v1, a13v2);
comparator c177 (a11v3, a13v4, a12v3, a14v4);
comparator c178 (a14v5, a13v6, a15v5, a14v6);
comparator c179 (a11v7, a12v8, a12v7, a13v8);
comparator c180 (a14v9, a15v10, a15v9, a16v10);
comparator c181 (a14v11, a13v12, a15v11, a14v12);
comparator c182 (a14v13, a12v14, a15v13, a13v14);
comparator c183 (a9v15, a9v16, a10v15, a10v16);
comparator c184 (a12v17, a14v18, a13v17, a15v18);
comparator c185 (a13v19, a14v20, a14v19, a15v20);
comparator c186 (a15v21, a14v22, a16v21, a15v22);
comparator c187 (a12v23, a11v24, a13v23, a12v24);
comparator c188 (a13v25, a14v26, a14v25, a15v26);
comparator c189 (a13v27, a11v28, a14v27, a12v28);
comparator c190 (a12v29, a9v30, a13v29, a10v30);
comparator c191 (a1v32, a1v33, a2v32, a2v33);
comparator c192 (a1v34, a1v35, a2v34, a2v35);
comparator c193 (a2v32, a2v34, a3v32, a3v34);
comparator c194 (a2v33, a2v35, a3v33, a3v35);
comparator c195 (a3v33, a3v34, a4v33, a4v34);
comparator c196 (a1v36, a1v37, a2v36, a2v37);
comparator c197 (a1v38, a1v39, a2v38, a2v39);
comparator c198 (a2v36, a2v38, a3v36, a3v38);
comparator c199 (a2v37, a2v39, a3v37, a3v39);
comparator c200 (a3v37, a3v38, a4v37, a4v38);
comparator c201 (a3v32, a3v36, a4v32, a4v36);
comparator c202 (a4v34, a4v38, a5v34, a5v38);
comparator c203 (a5v34, a4v36, a6v34, a5v36);
comparator c204 (a4v33, a4v37, a5v33, a5v37);
comparator c205 (a3v35, a3v39, a4v35, a4v39);
comparator c206 (a4v35, a5v37, a5v35, a6v37);
comparator c207 (a5v33, a6v34, a6v33, a7v34);
comparator c208 (a5v35, a5v36, a6v35, a6v36);
comparator c209 (a6v37, a5v38, a7v37, a6v38);
comparator c210 (a1v40, a1v41, a2v40, a2v41);
comparator c211 (a1v42, a1v43, a2v42, a2v43);
comparator c212 (a2v40, a2v42, a3v40, a3v42);
comparator c213 (a2v41, a2v43, a3v41, a3v43);
comparator c214 (a3v41, a3v42, a4v41, a4v42);
comparator c215 (a1v44, a1v45, a2v44, a2v45);
comparator c216 (a1v46, a1v47, a2v46, a2v47);
comparator c217 (a2v44, a2v46, a3v44, a3v46);
comparator c218 (a2v45, a2v47, a3v45, a3v47);
comparator c219 (a3v45, a3v46, a4v45, a4v46);
comparator c220 (a3v40, a3v44, a4v40, a4v44);
comparator c221 (a4v42, a4v46, a5v42, a5v46);
comparator c222 (a5v42, a4v44, a6v42, a5v44);
comparator c223 (a4v41, a4v45, a5v41, a5v45);
comparator c224 (a3v43, a3v47, a4v43, a4v47);
comparator c225 (a4v43, a5v45, a5v43, a6v45);
comparator c226 (a5v41, a6v42, a6v41, a7v42);
comparator c227 (a5v43, a5v44, a6v43, a6v44);
comparator c228 (a6v45, a5v46, a7v45, a6v46);
comparator c229 (a4v32, a4v40, a5v32, a5v40);
comparator c230 (a6v36, a6v44, a7v36, a7v44);
comparator c231 (a7v36, a5v40, a8v36, a6v40);
comparator c232 (a7v34, a7v42, a8v34, a8v42);
comparator c233 (a6v38, a6v46, a7v38, a7v46);
comparator c234 (a7v38, a8v42, a8v38, a9v42);
comparator c235 (a8v34, a8v36, a9v34, a9v36);
comparator c236 (a8v38, a6v40, a9v38, a7v40);
comparator c237 (a9v42, a7v44, a10v42, a8v44);
comparator c238 (a6v33, a6v41, a7v33, a7v41);
comparator c239 (a7v37, a7v45, a8v37, a8v45);
comparator c240 (a8v37, a7v41, a9v37, a8v41);
comparator c241 (a6v35, a6v43, a7v35, a7v43);
comparator c242 (a4v39, a4v47, a5v39, a5v47);
comparator c243 (a5v39, a7v43, a6v39, a8v43);
comparator c244 (a7v35, a9v37, a8v35, a10v37);
comparator c245 (a6v39, a8v41, a7v39, a9v41);
comparator c246 (a8v43, a8v45, a9v43, a9v45);
comparator c247 (a7v33, a9v34, a8v33, a10v34);
comparator c248 (a8v35, a9v36, a9v35, a10v36);
comparator c249 (a10v37, a9v38, a11v37, a10v38);
comparator c250 (a7v39, a7v40, a8v39, a8v40);
comparator c251 (a9v41, a10v42, a10v41, a11v42);
comparator c252 (a9v43, a8v44, a10v43, a9v44);
comparator c253 (a9v45, a7v46, a10v45, a8v46);
comparator c254 (a1v48, a1v49, a2v48, a2v49);
comparator c255 (a1v50, a1v51, a2v50, a2v51);
comparator c256 (a2v48, a2v50, a3v48, a3v50);
comparator c257 (a2v49, a2v51, a3v49, a3v51);
comparator c258 (a3v49, a3v50, a4v49, a4v50);
comparator c259 (a1v52, a1v53, a2v52, a2v53);
comparator c260 (a1v54, a1v55, a2v54, a2v55);
comparator c261 (a2v52, a2v54, a3v52, a3v54);
comparator c262 (a2v53, a2v55, a3v53, a3v55);
comparator c263 (a3v53, a3v54, a4v53, a4v54);
comparator c264 (a3v48, a3v52, a4v48, a4v52);
comparator c265 (a4v50, a4v54, a5v50, a5v54);
comparator c266 (a5v50, a4v52, a6v50, a5v52);
comparator c267 (a4v49, a4v53, a5v49, a5v53);
comparator c268 (a3v51, a3v55, a4v51, a4v55);
comparator c269 (a4v51, a5v53, a5v51, a6v53);
comparator c270 (a5v49, a6v50, a6v49, a7v50);
comparator c271 (a5v51, a5v52, a6v51, a6v52);
comparator c272 (a6v53, a5v54, a7v53, a6v54);
comparator c273 (a1v56, a1v57, a2v56, a2v57);
comparator c274 (a1v58, a1v59, a2v58, a2v59);
comparator c275 (a2v56, a2v58, a3v56, a3v58);
comparator c276 (a2v57, a2v59, a3v57, a3v59);
comparator c277 (a3v57, a3v58, a4v57, a4v58);
comparator c278 (a1v60, a1v61, a2v60, a2v61);
comparator c279 (a1v62, a1v63, a2v62, a2v63);
comparator c280 (a2v60, a2v62, a3v60, a3v62);
comparator c281 (a2v61, a2v63, a3v61, a3v63);
comparator c282 (a3v61, a3v62, a4v61, a4v62);
comparator c283 (a3v56, a3v60, a4v56, a4v60);
comparator c284 (a4v58, a4v62, a5v58, a5v62);
comparator c285 (a5v58, a4v60, a6v58, a5v60);
comparator c286 (a4v57, a4v61, a5v57, a5v61);
comparator c287 (a3v59, a3v63, a4v59, a4v63);
comparator c288 (a4v59, a5v61, a5v59, a6v61);
comparator c289 (a5v57, a6v58, a6v57, a7v58);
comparator c290 (a5v59, a5v60, a6v59, a6v60);
comparator c291 (a6v61, a5v62, a7v61, a6v62);
comparator c292 (a4v48, a4v56, a5v48, a5v56);
comparator c293 (a6v52, a6v60, a7v52, a7v60);
comparator c294 (a7v52, a5v56, a8v52, a6v56);
comparator c295 (a7v50, a7v58, a8v50, a8v58);
comparator c296 (a6v54, a6v62, a7v54, a7v62);
comparator c297 (a7v54, a8v58, a8v54, a9v58);
comparator c298 (a8v50, a8v52, a9v50, a9v52);
comparator c299 (a8v54, a6v56, a9v54, a7v56);
comparator c300 (a9v58, a7v60, a10v58, a8v60);
comparator c301 (a6v49, a6v57, a7v49, a7v57);
comparator c302 (a7v53, a7v61, a8v53, a8v61);
comparator c303 (a8v53, a7v57, a9v53, a8v57);
comparator c304 (a6v51, a6v59, a7v51, a7v59);
comparator c305 (a4v55, a4v63, a5v55, a5v63);
comparator c306 (a5v55, a7v59, a6v55, a8v59);
comparator c307 (a7v51, a9v53, a8v51, a10v53);
comparator c308 (a6v55, a8v57, a7v55, a9v57);
comparator c309 (a8v59, a8v61, a9v59, a9v61);
comparator c310 (a7v49, a9v50, a8v49, a10v50);
comparator c311 (a8v51, a9v52, a9v51, a10v52);
comparator c312 (a10v53, a9v54, a11v53, a10v54);
comparator c313 (a7v55, a7v56, a8v55, a8v56);
comparator c314 (a9v57, a10v58, a10v57, a11v58);
comparator c315 (a9v59, a8v60, a10v59, a9v60);
comparator c316 (a9v61, a7v62, a10v61, a8v62);
comparator c317 (a5v32, a5v48, a6v32, a6v48);
comparator c318 (a8v40, a8v56, a9v40, a9v56);
comparator c319 (a9v40, a6v48, a10v40, a7v48);
comparator c320 (a10v36, a10v52, a11v36, a11v52);
comparator c321 (a9v44, a9v60, a10v44, a10v60);
comparator c322 (a10v44, a11v52, a11v44, a12v52);
comparator c323 (a11v36, a10v40, a12v36, a11v40);
comparator c324 (a11v44, a7v48, a12v44, a8v48);
comparator c325 (a12v52, a9v56, a13v52, a10v56);
comparator c326 (a10v34, a10v50, a11v34, a11v50);
comparator c327 (a11v42, a11v58, a12v42, a12v58);
comparator c328 (a12v42, a11v50, a13v42, a12v50);
comparator c329 (a10v38, a10v54, a11v38, a11v54);
comparator c330 (a8v46, a8v62, a9v46, a9v62);
comparator c331 (a9v46, a11v54, a10v46, a12v54);
comparator c332 (a11v38, a13v42, a12v38, a14v42);
comparator c333 (a10v46, a12v50, a11v46, a13v50);
comparator c334 (a12v54, a12v58, a13v54, a13v58);
comparator c335 (a11v34, a12v36, a12v34, a13v36);
comparator c336 (a12v38, a11v40, a13v38, a12v40);
comparator c337 (a14v42, a12v44, a15v42, a13v44);
comparator c338 (a11v46, a8v48, a12v46, a9v48);
comparator c339 (a13v50, a13v52, a14v50, a14v52);
comparator c340 (a13v54, a10v56, a14v54, a11v56);
comparator c341 (a13v58, a10v60, a14v58, a11v60);
comparator c342 (a8v33, a8v49, a9v33, a9v49);
comparator c343 (a10v41, a10v57, a11v41, a11v57);
comparator c344 (a11v41, a9v49, a12v41, a10v49);
comparator c345 (a11v37, a11v53, a12v37, a12v53);
comparator c346 (a10v45, a10v61, a11v45, a11v61);
comparator c347 (a11v45, a12v53, a12v45, a13v53);
comparator c348 (a12v37, a12v41, a13v37, a13v41);
comparator c349 (a12v45, a10v49, a13v45, a11v49);
comparator c350 (a13v53, a11v57, a14v53, a12v57);
comparator c351 (a9v35, a9v51, a10v35, a10v51);
comparator c352 (a10v43, a10v59, a11v43, a11v59);
comparator c353 (a11v43, a10v51, a12v43, a11v51);
comparator c354 (a8v39, a8v55, a9v39, a9v55);
comparator c355 (a5v47, a5v63, a6v47, a6v63);
comparator c356 (a6v47, a9v55, a7v47, a10v55);
comparator c357 (a9v39, a12v43, a10v39, a13v43);
comparator c358 (a7v47, a11v51, a8v47, a12v51);
comparator c359 (a10v55, a11v59, a11v55, a12v59);
comparator c360 (a10v35, a13v37, a11v35, a14v37);
comparator c361 (a10v39, a13v41, a11v39, a14v41);
comparator c362 (a13v43, a13v45, a14v43, a14v45);
comparator c363 (a8v47, a11v49, a9v47, a12v49);
comparator c364 (a12v51, a14v53, a13v51, a15v53);
comparator c365 (a11v55, a12v57, a12v55, a13v57);
comparator c366 (a12v59, a11v61, a13v59, a12v61);
comparator c367 (a9v33, a12v34, a10v33, a13v34);
comparator c368 (a11v35, a13v36, a12v35, a14v36);
comparator c369 (a14v37, a13v38, a15v37, a14v38);
comparator c370 (a11v39, a12v40, a12v39, a13v40);
comparator c371 (a14v41, a15v42, a15v41, a16v42);
comparator c372 (a14v43, a13v44, a15v43, a14v44);
comparator c373 (a14v45, a12v46, a15v45, a13v46);
comparator c374 (a9v47, a9v48, a10v47, a10v48);
comparator c375 (a12v49, a14v50, a13v49, a15v50);
comparator c376 (a13v51, a14v52, a14v51, a15v52);
comparator c377 (a15v53, a14v54, a16v53, a15v54);
comparator c378 (a12v55, a11v56, a13v55, a12v56);
comparator c379 (a13v57, a14v58, a14v57, a15v58);
comparator c380 (a13v59, a11v60, a14v59, a12v60);
comparator c381 (a12v61, a9v62, a13v61, a10v62);
comparator c382 (a6v0, a6v32, a7v0, a7v32);
comparator c383 (a10v16, a10v48, a11v16, a11v48);
comparator c384 (a11v16, a7v32, a12v16, a8v32);
comparator c385 (a13v8, a13v40, a14v8, a14v40);
comparator c386 (a12v24, a12v56, a13v24, a13v56);
comparator c387 (a13v24, a14v40, a14v24, a15v40);
comparator c388 (a14v8, a12v16, a15v8, a13v16);
comparator c389 (a14v24, a8v32, a15v24, a9v32);
comparator c390 (a15v40, a11v48, a16v40, a12v48);
comparator c391 (a14v4, a14v36, a15v4, a15v36);
comparator c392 (a15v20, a15v52, a16v20, a16v52);
comparator c393 (a16v20, a15v36, a17v20, a16v36);
comparator c394 (a14v12, a14v44, a15v12, a15v44);
comparator c395 (a12v28, a12v60, a13v28, a13v60);
comparator c396 (a13v28, a15v44, a14v28, a16v44);
comparator c397 (a15v12, a17v20, a16v12, a18v20);
comparator c398 (a14v28, a16v36, a15v28, a17v36);
comparator c399 (a16v44, a16v52, a17v44, a17v52);
comparator c400 (a15v4, a15v8, a16v4, a16v8);
comparator c401 (a16v12, a13v16, a17v12, a14v16);
comparator c402 (a18v20, a15v24, a19v20, a16v24);
comparator c403 (a15v28, a9v32, a16v28, a10v32);
comparator c404 (a17v36, a16v40, a18v36, a17v40);
comparator c405 (a17v44, a12v48, a18v44, a13v48);
comparator c406 (a17v52, a13v56, a18v52, a14v56);
comparator c407 (a13v2, a13v34, a14v2, a14v34);
comparator c408 (a15v18, a15v50, a16v18, a16v50);
comparator c409 (a16v18, a14v34, a17v18, a15v34);
comparator c410 (a16v10, a16v42, a17v10, a17v42);
comparator c411 (a15v26, a15v58, a16v26, a16v58);
comparator c412 (a16v26, a17v42, a17v26, a18v42);
comparator c413 (a17v10, a17v18, a18v10, a18v18);
comparator c414 (a17v26, a15v34, a18v26, a16v34);
comparator c415 (a18v42, a16v50, a19v42, a17v50);
comparator c416 (a14v6, a14v38, a15v6, a15v38);
comparator c417 (a15v22, a15v54, a16v22, a16v54);
comparator c418 (a16v22, a15v38, a17v22, a16v38);
comparator c419 (a13v14, a13v46, a14v14, a14v46);
comparator c420 (a10v30, a10v62, a11v30, a11v62);
comparator c421 (a11v30, a14v46, a12v30, a15v46);
comparator c422 (a14v14, a17v22, a15v14, a18v22);
comparator c423 (a12v30, a16v38, a13v30, a17v38);
comparator c424 (a15v46, a16v54, a16v46, a17v54);
comparator c425 (a15v6, a18v10, a16v6, a19v10);
comparator c426 (a15v14, a18v18, a16v14, a19v18);
comparator c427 (a18v22, a18v26, a19v22, a19v26);
comparator c428 (a13v30, a16v34, a14v30, a17v34);
comparator c429 (a17v38, a19v42, a18v38, a20v42);
comparator c430 (a16v46, a17v50, a17v46, a18v50);
comparator c431 (a17v54, a16v58, a18v54, a17v58);
comparator c432 (a14v2, a16v4, a15v2, a17v4);
comparator c433 (a16v6, a16v8, a17v6, a17v8);
comparator c434 (a19v10, a17v12, a20v10, a18v12);
comparator c435 (a16v14, a14v16, a17v14, a15v16);
comparator c436 (a19v18, a19v20, a20v18, a20v20);
comparator c437 (a19v22, a16v24, a20v22, a17v24);
comparator c438 (a19v26, a16v28, a20v26, a17v28);
comparator c439 (a14v30, a10v32, a15v30, a11v32);
comparator c440 (a17v34, a18v36, a18v34, a19v36);
comparator c441 (a18v38, a17v40, a19v38, a18v40);
comparator c442 (a20v42, a18v44, a21v42, a19v44);
comparator c443 (a17v46, a13v48, a18v46, a14v48);
comparator c444 (a18v50, a18v52, a19v50, a19v52);
comparator c445 (a18v54, a14v56, a19v54, a15v56);
comparator c446 (a17v58, a13v60, a18v58, a14v60);
comparator c447 (a10v1, a10v33, a11v1, a11v33);
comparator c448 (a13v17, a13v49, a14v17, a14v49);
comparator c449 (a14v17, a11v33, a15v17, a12v33);
comparator c450 (a15v9, a15v41, a16v9, a16v41);
comparator c451 (a14v25, a14v57, a15v25, a15v57);
comparator c452 (a15v25, a16v41, a16v25, a17v41);
comparator c453 (a16v9, a15v17, a17v9, a16v17);
comparator c454 (a16v25, a12v33, a17v25, a13v33);
comparator c455 (a17v41, a14v49, a18v41, a15v49);
comparator c456 (a15v5, a15v37, a16v5, a16v37);
comparator c457 (a16v21, a16v53, a17v21, a17v53);
comparator c458 (a17v21, a16v37, a18v21, a17v37);
comparator c459 (a15v13, a15v45, a16v13, a16v45);
comparator c460 (a13v29, a13v61, a14v29, a14v61);
comparator c461 (a14v29, a16v45, a15v29, a17v45);
comparator c462 (a16v13, a18v21, a17v13, a19v21);
comparator c463 (a15v29, a17v37, a16v29, a18v37);
comparator c464 (a17v45, a17v53, a18v45, a18v53);
comparator c465 (a16v5, a17v9, a17v5, a18v9);
comparator c466 (a17v13, a16v17, a18v13, a17v17);
comparator c467 (a19v21, a17v25, a20v21, a18v25);
comparator c468 (a16v29, a13v33, a17v29, a14v33);
comparator c469 (a18v37, a18v41, a19v37, a19v41);
comparator c470 (a18v45, a15v49, a19v45, a16v49);
comparator c471 (a18v53, a15v57, a19v53, a16v57);
comparator c472 (a12v3, a12v35, a13v3, a13v35);
comparator c473 (a14v19, a14v51, a15v19, a15v51);
comparator c474 (a15v19, a13v35, a16v19, a14v35);
comparator c475 (a15v11, a15v43, a16v11, a16v43);
comparator c476 (a14v27, a14v59, a15v27, a15v59);
comparator c477 (a15v27, a16v43, a16v27, a17v43);
comparator c478 (a16v11, a16v19, a17v11, a17v19);
comparator c479 (a16v27, a14v35, a17v27, a15v35);
comparator c480 (a17v43, a15v51, a18v43, a16v51);
comparator c481 (a12v7, a12v39, a13v7, a13v39);
comparator c482 (a13v23, a13v55, a14v23, a14v55);
comparator c483 (a14v23, a13v39, a15v23, a14v39);
comparator c484 (a10v15, a10v47, a11v15, a11v47);
comparator c485 (a6v31, a6v63, a7v31, a7v63);
comparator c486 (a7v31, a11v47, a8v31, a12v47);
comparator c487 (a11v15, a15v23, a12v15, a16v23);
comparator c488 (a8v31, a14v39, a9v31, a15v39);
comparator c489 (a12v47, a14v55, a13v47, a15v55);
comparator c490 (a13v7, a17v11, a14v7, a18v11);
comparator c491 (a12v15, a17v19, a13v15, a18v19);
comparator c492 (a16v23, a17v27, a17v23, a18v27);
comparator c493 (a9v31, a15v35, a10v31, a16v35);
comparator c494 (a15v39, a18v43, a16v39, a19v43);
comparator c495 (a13v47, a16v51, a14v47, a17v51);
comparator c496 (a15v55, a15v59, a16v55, a16v59);
comparator c497 (a13v3, a17v5, a14v3, a18v5);
comparator c498 (a14v7, a18v9, a15v7, a19v9);
comparator c499 (a18v11, a18v13, a19v11, a19v13);
comparator c500 (a13v15, a17v17, a14v15, a18v17);
comparator c501 (a18v19, a20v21, a19v19, a21v21);
comparator c502 (a17v23, a18v25, a18v23, a19v25);
comparator c503 (a18v27, a17v29, a19v27, a18v29);
comparator c504 (a10v31, a14v33, a11v31, a15v33);
comparator c505 (a16v35, a19v37, a17v35, a20v37);
comparator c506 (a16v39, a19v41, a17v39, a20v41);
comparator c507 (a19v43, a19v45, a20v43, a20v45);
comparator c508 (a14v47, a16v49, a15v47, a17v49);
comparator c509 (a17v51, a19v53, a18v51, a20v53);
comparator c510 (a16v55, a16v57, a17v55, a17v57);
comparator c511 (a16v59, a14v61, a17v59, a15v61);
comparator c512 (a11v1, a15v2, a12v1, a16v2);
comparator c513 (a14v3, a17v4, a15v3, a18v4);
comparator c514 (a18v5, a17v6, a19v5, a18v6);
comparator c515 (a15v7, a17v8, a16v7, a18v8);
comparator c516 (a19v9, a20v10, a20v9, a21v10);
comparator c517 (a19v11, a18v12, a20v11, a19v12);
comparator c518 (a19v13, a17v14, a20v13, a18v14);
comparator c519 (a14v15, a15v16, a15v15, a16v16);
comparator c520 (a18v17, a20v18, a19v17, a21v18);
comparator c521 (a19v19, a20v20, a20v19, a21v20);
comparator c522 (a21v21, a20v22, a22v21, a21v22);
comparator c523 (a18v23, a17v24, a19v23, a18v24);
comparator c524 (a19v25, a20v26, a20v25, a21v26);
comparator c525 (a19v27, a17v28, a20v27, a18v28);
comparator c526 (a18v29, a15v30, a19v29, a16v30);
comparator c527 (a11v31, a11v32, a12v31, a12v32);
comparator c528 (a15v33, a18v34, a16v33, a19v34);
comparator c529 (a17v35, a19v36, a18v35, a20v36);
comparator c530 (a20v37, a19v38, a21v37, a20v38);
comparator c531 (a17v39, a18v40, a18v39, a19v40);
comparator c532 (a20v41, a21v42, a21v41, a22v42);
comparator c533 (a20v43, a19v44, a21v43, a20v44);
comparator c534 (a20v45, a18v46, a21v45, a19v46);
comparator c535 (a15v47, a14v48, a16v47, a15v48);
comparator c536 (a17v49, a19v50, a18v49, a20v50);
comparator c537 (a18v51, a19v52, a19v51, a20v52);
comparator c538 (a20v53, a19v54, a21v53, a20v54);
comparator c539 (a17v55, a15v56, a18v55, a16v56);
comparator c540 (a17v57, a18v58, a18v57, a19v58);
comparator c541 (a17v59, a14v60, a18v59, a15v60);
comparator c542 (a15v61, a11v62, a16v61, a12v62);


endmodule

module bsort_49(data_in, data_out);


input   [391:0] data_in;
output  [7:0] data_out;

wire    [511:0] c_in;
wire    [511:0] c_out;

assign  c_in[391:0]   = data_in;
assign  c_in[511:392] = 0;

assign  data_out[3:0] = c_out[315:312];
assign  data_out[7:4] = c_out[319:316];
bsort b1(.data_in(c_in), .data_out(c_out));


endmodule
module LMFE ( clk, reset, Din, in_en, busy, out_valid, Dout);
input          clk;
input          reset;
input          in_en;
output         busy;
output         out_valid;
input   [7:0]  Din;
output  [7:0]  Dout;

integer i;

parameter STATUS_IDLE  = 2'b00
        , STATUS_WRITE = 2'b11
        , STATUS_READ  = 2'b10;

reg [7:0] Din_2;
always @ (posedge clk) begin
    Din_2 <= (reset) ? 0 : Din;
end


reg [55:0] filter1; // 8bits x 7 pixels
reg [55:0] filter2;
reg [55:0] filter3;
reg [55:0] filter4;
reg [55:0] filter5;
reg [55:0] filter6;
reg [55:0] filter;

reg  [3:0] in_ctrl   [8:0];

wire [7:0]  sram_out      [8:0]; // 1+7, 0:   zonst_zero
reg  [1:0]  s_ctrl        [8:0]; // For 8 sram, sram_overall_ctrl
                         // 0: null, 1:8: sram
assign sram_out[0] = 0;


// TODO: NOTE sram_en only slow 1 clock, while data in slow 2 clock
sram_ctrl sram1(.clk(clk), .reset(reset), .sram_in_ctrl(s_ctrl[1])
                     , .sram_in(Din_2), .sram_out(sram_out[1]));
sram_ctrl sram2(.clk(clk), .reset(reset), .sram_in_ctrl(s_ctrl[2])
                     , .sram_in(Din_2), .sram_out(sram_out[2]));
sram_ctrl sram3(.clk(clk), .reset(reset), .sram_in_ctrl(s_ctrl[3])
                     , .sram_in(Din_2), .sram_out(sram_out[3]));
sram_ctrl sram4(.clk(clk), .reset(reset), .sram_in_ctrl(s_ctrl[4])
                      , .sram_in(Din_2), .sram_out(sram_out[4]));
sram_ctrl sram5(.clk(clk), .reset(reset), .sram_in_ctrl(s_ctrl[5])
                     , .sram_in(Din_2), .sram_out(sram_out[5]));
sram_ctrl sram6(.clk(clk), .reset(reset), .sram_in_ctrl(s_ctrl[6])
                     , .sram_in(Din_2), .sram_out(sram_out[6]));
sram_ctrl sram7(.clk(clk), .reset(reset), .sram_in_ctrl(s_ctrl[7])
                     , .sram_in(Din_2), .sram_out(sram_out[7]));
sram_ctrl sram8(.clk(clk), .reset(reset), .sram_in_ctrl(s_ctrl[8])
                     , .sram_in(Din_2), .sram_out(sram_out[8]));


reg [7:0] filter_in [6:0];

reg [7:0] counter_seq;

always @ (posedge clk) begin
    for(i = 0; i<7; i = i+1)
        filter_in[i] <= sram_out[in_ctrl[i]];
end
// filter1 ... filter6 filter <= sram_data
always @ (posedge clk) begin
    if(reset) begin
        filter1 <= 0;
        filter2 <= 0;
        filter3 <= 0;
        filter4 <= 0;
        filter5 <= 0;
        filter6 <= 0;
        filter <= 0;
    end
    else begin
    filter1 <= filter2;
    filter2 <= filter3;
    filter3 <= filter4;
    filter4 <= filter5;
    filter5 <= filter6;
    filter6 <= filter;
    filter  <= (counter_seq == 8'h00 || counter_seq == 8'h01 || counter_seq == 8'h02)  // test
             ? 0 
             : {filter_in[0], filter_in[1], filter_in[2]
    , filter_in[3], filter_in[4], filter_in[5], filter_in[6]};
    end
end

wire  [391:0] sort_in;
wire  [7:0]   sort_out;

bsort_49 b1(.data_in(sort_in), .data_out(sort_out));
assign sort_in = { filter1, filter2, filter3, filter4
                 , filter5, filter6, filter};
assign Dout = sort_out;

reg  [2:0]  state;
reg  [2:0]  next_state;

reg [1:0] seq_read;
reg [1:0] seq_write;
reg [1:0] seq_idle;
assign busy = (counter_seq < 3) ? 1'b1 : 1'b0;
always @ (posedge clk) begin
    seq_idle <= STATUS_IDLE;
    if(reset) begin
        seq_write <= STATUS_IDLE;
        seq_read <= STATUS_IDLE;
    end
    else begin
        seq_write <= (counter_seq < 3) ? STATUS_IDLE : STATUS_WRITE;
        seq_read  <= (counter_seq < 3) ? STATUS_IDLE : STATUS_READ;
    end
end
always @ (posedge clk) begin
    if(reset) begin
        counter_seq <= 0;
    end
    else begin
        counter_seq <= (counter_seq == 130) ? 0 : counter_seq + 1'b1;
    end
end


reg  [7:0] state_select;
reg  [1:0] select [8:0];
wire all_clk;
parameter WW  = 2'b11    // write
        , WR  = 2'b10   // read 
        , WI  = 2'b00;  // idle
parameter INS0 = 4'b0000
        , INS1 = INS0 + 1'b1
        , INS2 = INS1 + 1'b1
        , INS3 = INS2 + 1'b1
        , INS4 = INS3 + 1'b1
        , INS5 = INS4 + 1'b1
        , INS6 = INS5 + 1'b1
        , INS7 = INS6 + 1'b1
        , INS8 = INS7 + 1'b1;
               // 8   7   6   5   4   3   2   1   0
parameter W1  =  {WI, WI, WI, WI, WI, WI, WI, WW, WI};
parameter W2  =  {WI, WI, WI, WW, WR, WR, WR, WR, WI};
parameter II  =  {INS0,INS0,INS0,INS0,INS0,INS0,INS0,INS0};
parameter I1  =  {INS5,INS4,INS3,INS2,INS1,INS0,INS0,INS0};
parameter I2  =  {INS6,INS5,INS4,INS3,INS2,INS1,INS0,INS0};
parameter I3  =  {INS7,INS6,INS5,INS4,INS3,INS2,INS1,INS0};
parameter I4  =  {INS8,INS7,INS6,INS5,INS4,INS3,INS2,INS1};
reg [17:0]  to_w_r;
reg [31:0]  to_ctrl;

always @ (posedge all_clk) begin
    if(reset)
        to_ctrl <= II;
    else begin
        case(state_select)
            8'h03: to_ctrl <= I1;
            8'h04: to_ctrl <= I2;
            8'h05: to_ctrl <= I3;
            8'h06: to_ctrl <= I4;
            8'h7f: to_ctrl <= { INS0, to_ctrl[31:4] };
            8'h80: to_ctrl <= { INS0, to_ctrl[31:4] };
            8'h81: to_ctrl <= { INS0, to_ctrl[31:4] };
            8'h82: to_ctrl <= { INS0, to_ctrl[31:4] };
            default: to_ctrl <= { to_ctrl[3:0], to_ctrl[31:4]};
        endcase
    end
end
always @ (posedge all_clk) begin
    if(reset)
        to_w_r <= W1;
    else begin
        case(state_select)
            7'h03: to_w_r         <= W2; // 4-1
            7'h04: to_w_r[17:2]   <= (to_w_r[17:2] << 2)+WR;
            7'h05: to_w_r[17:2]   <= (to_w_r[17:2] << 2)+WR;
            7'h06: to_w_r[17:2]   <= (to_w_r[17:2] << 2)+WR;
            8'h80: to_w_r[17:2]   <= (to_w_r[17:2] << 2)+WI;
            8'h81: to_w_r[17:2]   <= (to_w_r[17:2] << 2)+WI;
            8'h82: to_w_r[17:2]   <= (to_w_r[17:2] << 2)+WI;
            default: to_w_r[17:2] <= { to_w_r[15:2], to_w_r[17:16] };
        endcase
    end
end

always @ (*) begin
    case(state_select)
        default: begin
            { select[8], select[7], select[6], select[5]
            , select[4], select[3], select[2], select[1], select[0] } = to_w_r;
            { in_ctrl[6], in_ctrl[5], in_ctrl[4], in_ctrl[3]
            , in_ctrl[2], in_ctrl[1], in_ctrl[0] } = to_ctrl;
        end
    endcase
end


always @ (posedge all_clk) begin
    if(reset) begin
        state_select <= 0;
    end
    else begin
        state_select <= state_select+1'b1; // TODO: determine length
    end
end

always @ (*) begin
    for(i=0; i<9; i = i+1)
        s_ctrl[i] = select[i];
end

assign all_clk = (seq_read == STATUS_IDLE) ? 1'b1 : 1'b0;


reg out_valid_reg;
reg o1, o2, o3;
always @ (posedge clk) begin
    o1 <= !busy;
    o2 <= o1;
    o3 <= o2;
end
always @ (posedge clk) begin
    if(reset) out_valid_reg <= 1'b0;
    else begin
    if(state_select > 3)
        if(state_select == 4)
            out_valid_reg <= (counter_seq > 5 || counter_seq ==0) ? 1'b1 : 1'b0;
        else
            out_valid_reg <= o3;
    end
end
assign out_valid = out_valid_reg;

endmodule
