module mem(clk);

reg [3:0] mem_array [2:0];

endmodule
