module A(reset);
input reset;
parameter PARA_A = 10;
endmodule
